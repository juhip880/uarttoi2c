jangnkl
